`timescale 1ns / 1ps

module ALU(
	input [31:0]a,
	input [31:0]b,
	input [2:0]alucont,
	output reg [31:0]result,
	output zero
);

reg sltresult=0;
always @(*)
    begin
    if(a[31] == b[31]) sltresult = (a<b);
    else if(a[31]==1) sltresult = 1;
    else sltresult = 0;  
    end

always @(*)
case(alucont)
3'b000: result = a&b; //and
3'b001: result = a|b; //or
3'b010: result = a+b; //add
3'b011: result = b << a; //not used
3'b100: result = b[31]==0?(b>>a):((b >> a) | ( ( (32'b11111111111111111111111111111111) >> (32-a)  ) << (32-a) ));//SRA
3'b101: result = b >> a;//SRL
3'b110: result = a-b; //sub
3'b111: result = sltresult;//slt
endcase

assign #1 zero = !result;

endmodule


